library verilog;
use verilog.vl_types.all;
entity light_show is
    port(
        light_clk       : in     vl_logic;
        SW_choose       : in     vl_logic;
        check_in        : in     vl_logic_vector(7 downto 0);
        read            : in     vl_logic;
        write           : in     vl_logic;
        arload          : in     vl_logic;
        arinc           : in     vl_logic;
        pcinc           : in     vl_logic;
        pcload          : in     vl_logic;
        drload          : in     vl_logic;
        trload          : in     vl_logic;
        irload          : in     vl_logic;
        rload           : in     vl_logic;
        acload          : in     vl_logic;
        zload           : in     vl_logic;
        pcbus           : in     vl_logic;
        drhbus          : in     vl_logic_vector(15 downto 8);
        drlbus          : in     vl_logic_vector(7 downto 0);
        trbus           : in     vl_logic;
        rbus            : in     vl_logic;
        acbus           : in     vl_logic;
        membus          : in     vl_logic;
        busmem          : in     vl_logic;
        clr             : in     vl_logic;
        State           : in     vl_logic_vector(1 downto 0);
        MAR             : in     vl_logic_vector(7 downto 0);
        AC              : in     vl_logic_vector(7 downto 0);
        R               : in     vl_logic_vector(7 downto 0);
        Z               : in     vl_logic;
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        HEX4            : out    vl_logic_vector(6 downto 0);
        HEX5            : out    vl_logic_vector(6 downto 0);
        HEX6            : out    vl_logic_vector(6 downto 0);
        HEX7            : out    vl_logic_vector(6 downto 0);
        State_LED       : out    vl_logic_vector(1 downto 0);
        quick_low_led   : out    vl_logic;
        read_led        : in     vl_logic;
        write_led       : in     vl_logic;
        arload_led      : in     vl_logic;
        arinc_led       : in     vl_logic;
        pcinc_led       : in     vl_logic;
        pcload_led      : in     vl_logic;
        drload_led      : in     vl_logic;
        trload_led      : in     vl_logic;
        irload_led      : in     vl_logic;
        rload_led       : in     vl_logic;
        acload_led      : in     vl_logic;
        zload_led       : in     vl_logic;
        pcbus_led       : in     vl_logic;
        drhbus_led      : in     vl_logic;
        drlbus_led      : in     vl_logic;
        trbus_led       : in     vl_logic;
        rbus_led        : in     vl_logic;
        acbus_led       : in     vl_logic;
        membus_led      : in     vl_logic;
        busmem_led      : in     vl_logic;
        clr_led         : in     vl_logic
    );
end light_show;
